module decoder (
input reg[]
);

